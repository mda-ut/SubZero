// DE0_Nano_SOPC.v

// Generated using ACDS version 13.1 162 at 2015.07.25.01:54:10

`timescale 1 ps / 1 ps
module DE0_Nano_SOPC (
		input  wire        reset_n,                                   //                  clk_50_clk_in_reset.reset_n
		input  wire        clk_50,                                    //                        clk_50_clk_in.clk
		input  wire [1:0]  in_port_to_the_key,                        //              key_external_connection.export
		input  wire [3:0]  in_port_to_the_sw,                         //               sw_external_connection.export
		output wire [7:0]  out_port_from_the_led,                     //              led_external_connection.export
		output wire        out_port_from_the_i2c_scl,                 //          i2c_scl_external_connection.export
		inout  wire        bidir_port_to_and_from_the_i2c_sda,        //          i2c_sda_external_connection.export
		output wire [12:0] zs_addr_from_the_sdram,                    //                           sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,                      //                                     .ba
		output wire        zs_cas_n_from_the_sdram,                   //                                     .cas_n
		output wire        zs_cke_from_the_sdram,                     //                                     .cke
		output wire        zs_cs_n_from_the_sdram,                    //                                     .cs_n
		inout  wire [15:0] zs_dq_to_and_from_the_sdram,               //                                     .dq
		output wire [1:0]  zs_dqm_from_the_sdram,                     //                                     .dqm
		output wire        zs_ras_n_from_the_sdram,                   //                                     .ras_n
		output wire        zs_we_n_from_the_sdram,                    //                                     .we_n
		output wire        altpll_sys,                                //                           c0_out_clk.clk
		output wire        altpll_sdram,                              //                        altpll_sys_c1.clk
		output wire        altpll_io,                                 //                           c2_out_clk.clk
		output wire        altpll_sys_c3_out,                         //                        altpll_sys_c3.clk
		output wire        altpll_adc,                                //                           c4_out_clk.clk
		output wire        locked_from_the_altpll_sys,                //            altpll_sys_locked_conduit.export
		output wire        phasedone_from_the_altpll_sys,             //         altpll_sys_phasedone_conduit.export
		input  wire        in_port_to_the_g_sensor_int,               //     g_sensor_int_external_connection.export
		output wire        dclk_from_the_epcs,                        //                        epcs_external.dclk
		output wire        sce_from_the_epcs,                         //                                     .sce
		output wire        sdo_from_the_epcs,                         //                                     .sdo
		input  wire        data0_to_the_epcs,                         //                                     .data0
		inout  wire        SPI_SDIO_to_and_from_the_gsensor_spi,      //              gsensor_spi_conduit_end.SDIO
		output wire        SPI_SCLK_from_the_gsensor_spi,             //                                     .SCLK
		output wire        SPI_CS_n_from_the_gsensor_spi,             //                                     .CS_n
		output wire        out_port_from_the_select_i2c_clk,          //   select_i2c_clk_external_connection.export
		output wire [23:0] GPIO_out_from_the_motor_controller_0,      //       motor_controller_0_conduit_end.export
		output wire        kill_sw_from_the_power_management_slave_0, // power_management_slave_0_conduit_end.kill_sw
		output wire [2:0]  mux_from_the_power_management_slave_0,     //                                     .mux
		input  wire        data_to_the_power_management_slave_0,      //                                     .data
		input  wire        sys_clk_to_the_imu_controller_0,           //         imu_controller_0_conduit_end.sys_clk
		input  wire        ADC_SDAT_to_the_imu_controller_0,          //                                     .ADC_SDAT
		output wire        ADC_CS_N_from_the_imu_controller_0,        //                                     .ADC_CS_N
		output wire        ADC_SADDR_from_the_imu_controller_0,       //                                     .ADC_SADDR
		output wire        ADC_SCLK_from_the_imu_controller_0,        //                                     .ADC_SCLK
		input  wire        UART_RXD_to_the_RS232_0,                   //                  RS232_0_conduit_end.export
		output wire        UART_TXD_from_the_RS232_0                  //                RS232_0_conduit_end_1.export
	);

	wire   [3:0] mm_interconnect_0_imu_controller_0_avalon_slave_0_address;            // mm_interconnect_0:imu_controller_0_avalon_slave_0_address -> imu_controller_0:addr
	wire         mm_interconnect_0_imu_controller_0_avalon_slave_0_chipselect;         // mm_interconnect_0:imu_controller_0_avalon_slave_0_chipselect -> imu_controller_0:chipselect
	wire         mm_interconnect_0_imu_controller_0_avalon_slave_0_read;               // mm_interconnect_0:imu_controller_0_avalon_slave_0_read -> imu_controller_0:read
	wire  [31:0] mm_interconnect_0_imu_controller_0_avalon_slave_0_readdata;           // imu_controller_0:readdata -> mm_interconnect_0:imu_controller_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_clock_crossing_io2_s0_waitrequest;                  // clock_crossing_io2:s0_waitrequest -> mm_interconnect_0:clock_crossing_io2_s0_waitrequest
	wire   [0:0] mm_interconnect_0_clock_crossing_io2_s0_burstcount;                   // mm_interconnect_0:clock_crossing_io2_s0_burstcount -> clock_crossing_io2:s0_burstcount
	wire  [31:0] mm_interconnect_0_clock_crossing_io2_s0_writedata;                    // mm_interconnect_0:clock_crossing_io2_s0_writedata -> clock_crossing_io2:s0_writedata
	wire  [11:0] mm_interconnect_0_clock_crossing_io2_s0_address;                      // mm_interconnect_0:clock_crossing_io2_s0_address -> clock_crossing_io2:s0_address
	wire         mm_interconnect_0_clock_crossing_io2_s0_write;                        // mm_interconnect_0:clock_crossing_io2_s0_write -> clock_crossing_io2:s0_write
	wire         mm_interconnect_0_clock_crossing_io2_s0_read;                         // mm_interconnect_0:clock_crossing_io2_s0_read -> clock_crossing_io2:s0_read
	wire  [31:0] mm_interconnect_0_clock_crossing_io2_s0_readdata;                     // clock_crossing_io2:s0_readdata -> mm_interconnect_0:clock_crossing_io2_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io2_s0_debugaccess;                  // mm_interconnect_0:clock_crossing_io2_s0_debugaccess -> clock_crossing_io2:s0_debugaccess
	wire         mm_interconnect_0_clock_crossing_io2_s0_readdatavalid;                // clock_crossing_io2:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io2_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_clock_crossing_io2_s0_byteenable;                   // mm_interconnect_0:clock_crossing_io2_s0_byteenable -> clock_crossing_io2:s0_byteenable
	wire  [15:0] mm_interconnect_0_controller_interrupt_counter_s1_writedata;          // mm_interconnect_0:controller_interrupt_counter_s1_writedata -> controller_interrupt_counter:writedata
	wire   [2:0] mm_interconnect_0_controller_interrupt_counter_s1_address;            // mm_interconnect_0:controller_interrupt_counter_s1_address -> controller_interrupt_counter:address
	wire         mm_interconnect_0_controller_interrupt_counter_s1_chipselect;         // mm_interconnect_0:controller_interrupt_counter_s1_chipselect -> controller_interrupt_counter:chipselect
	wire         mm_interconnect_0_controller_interrupt_counter_s1_write;              // mm_interconnect_0:controller_interrupt_counter_s1_write -> controller_interrupt_counter:write_n
	wire  [15:0] mm_interconnect_0_controller_interrupt_counter_s1_readdata;           // controller_interrupt_counter:readdata -> mm_interconnect_0:controller_interrupt_counter_s1_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;            // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;               // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                  // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                    // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                      // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                        // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                         // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                     // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                  // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                   // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;                   // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;                    // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;                     // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire   [6:0] mm_interconnect_0_clock_crossing_io_s0_address;                       // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_write;                         // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire         mm_interconnect_0_clock_crossing_io_s0_read;                          // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;                      // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;                   // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;                 // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;                    // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         cpu_data_master_waitrequest;                                          // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                            // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [26:0] cpu_data_master_address;                                              // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                                // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                                 // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                             // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                          // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                           // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_instruction_master_waitrequest;                                   // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                                       // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                          // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                      // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire  [31:0] mm_interconnect_0_power_management_slave_0_avalon_slave_0_writedata;  // mm_interconnect_0:power_management_slave_0_avalon_slave_0_writedata -> power_management_slave_0:writedata
	wire         mm_interconnect_0_power_management_slave_0_avalon_slave_0_chipselect; // mm_interconnect_0:power_management_slave_0_avalon_slave_0_chipselect -> power_management_slave_0:chipselect
	wire         mm_interconnect_0_power_management_slave_0_avalon_slave_0_write;      // mm_interconnect_0:power_management_slave_0_avalon_slave_0_write -> power_management_slave_0:write
	wire         mm_interconnect_0_power_management_slave_0_avalon_slave_0_read;       // mm_interconnect_0:power_management_slave_0_avalon_slave_0_read -> power_management_slave_0:read
	wire  [31:0] mm_interconnect_0_power_management_slave_0_avalon_slave_0_readdata;   // power_management_slave_0:readdata -> mm_interconnect_0:power_management_slave_0_avalon_slave_0_readdata
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_writedata;                     // mm_interconnect_0:altpll_sys_pll_slave_writedata -> altpll_sys:writedata
	wire   [1:0] mm_interconnect_0_altpll_sys_pll_slave_address;                       // mm_interconnect_0:altpll_sys_pll_slave_address -> altpll_sys:address
	wire         mm_interconnect_0_altpll_sys_pll_slave_write;                         // mm_interconnect_0:altpll_sys_pll_slave_write -> altpll_sys:write
	wire         mm_interconnect_0_altpll_sys_pll_slave_read;                          // mm_interconnect_0:altpll_sys_pll_slave_read -> altpll_sys:read
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_readdata;                      // altpll_sys:readdata -> mm_interconnect_0:altpll_sys_pll_slave_readdata
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_slave_0_writedata;                   // mm_interconnect_0:RS232_0_avalon_slave_0_writedata -> RS232_0:writedata
	wire   [0:0] mm_interconnect_0_rs232_0_avalon_slave_0_address;                     // mm_interconnect_0:RS232_0_avalon_slave_0_address -> RS232_0:address
	wire         mm_interconnect_0_rs232_0_avalon_slave_0_chipselect;                  // mm_interconnect_0:RS232_0_avalon_slave_0_chipselect -> RS232_0:chipselect
	wire         mm_interconnect_0_rs232_0_avalon_slave_0_write;                       // mm_interconnect_0:RS232_0_avalon_slave_0_write -> RS232_0:write
	wire         mm_interconnect_0_rs232_0_avalon_slave_0_read;                        // mm_interconnect_0:RS232_0_avalon_slave_0_read -> RS232_0:read
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_slave_0_readdata;                    // RS232_0:readdata -> mm_interconnect_0:RS232_0_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_0_rs232_0_avalon_slave_0_byteenable;                  // mm_interconnect_0:RS232_0_avalon_slave_0_byteenable -> RS232_0:byteenable
	wire         mm_interconnect_0_sdram_s1_waitrequest;                               // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                 // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                   // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                                // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                     // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                      // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                  // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                             // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [31:0] mm_interconnect_0_motor_controller_0_avalon_slave_0_writedata;        // mm_interconnect_0:motor_controller_0_avalon_slave_0_writedata -> motor_controller_0:writedata
	wire   [3:0] mm_interconnect_0_motor_controller_0_avalon_slave_0_address;          // mm_interconnect_0:motor_controller_0_avalon_slave_0_address -> motor_controller_0:addr
	wire         mm_interconnect_0_motor_controller_0_avalon_slave_0_chipselect;       // mm_interconnect_0:motor_controller_0_avalon_slave_0_chipselect -> motor_controller_0:chipselect
	wire         mm_interconnect_0_motor_controller_0_avalon_slave_0_write;            // mm_interconnect_0:motor_controller_0_avalon_slave_0_write -> motor_controller_0:write
	wire  [31:0] mm_interconnect_1_sw_s1_writedata;                                    // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                                      // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_sw_s1_chipselect;                                   // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire         mm_interconnect_1_sw_s1_write;                                        // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                                     // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                                   // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire   [1:0] mm_interconnect_1_key_s1_address;                                     // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_chipselect;                                  // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire         mm_interconnect_1_key_s1_write;                                       // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                                    // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                                   // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire   [1:0] mm_interconnect_1_led_s1_address;                                     // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_chipselect;                                  // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire         mm_interconnect_1_led_s1_write;                                       // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                                    // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire  [31:0] mm_interconnect_1_select_i2c_clk_s1_writedata;                        // mm_interconnect_1:select_i2c_clk_s1_writedata -> select_i2c_clk:writedata
	wire   [1:0] mm_interconnect_1_select_i2c_clk_s1_address;                          // mm_interconnect_1:select_i2c_clk_s1_address -> select_i2c_clk:address
	wire         mm_interconnect_1_select_i2c_clk_s1_chipselect;                       // mm_interconnect_1:select_i2c_clk_s1_chipselect -> select_i2c_clk:chipselect
	wire         mm_interconnect_1_select_i2c_clk_s1_write;                            // mm_interconnect_1:select_i2c_clk_s1_write -> select_i2c_clk:write_n
	wire  [31:0] mm_interconnect_1_select_i2c_clk_s1_readdata;                         // select_i2c_clk:readdata -> mm_interconnect_1:select_i2c_clk_s1_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                        // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                       // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire  [31:0] mm_interconnect_1_g_sensor_int_s1_writedata;                          // mm_interconnect_1:g_sensor_int_s1_writedata -> g_sensor_int:writedata
	wire   [1:0] mm_interconnect_1_g_sensor_int_s1_address;                            // mm_interconnect_1:g_sensor_int_s1_address -> g_sensor_int:address
	wire         mm_interconnect_1_g_sensor_int_s1_chipselect;                         // mm_interconnect_1:g_sensor_int_s1_chipselect -> g_sensor_int:chipselect
	wire         mm_interconnect_1_g_sensor_int_s1_write;                              // mm_interconnect_1:g_sensor_int_s1_write -> g_sensor_int:write_n
	wire  [31:0] mm_interconnect_1_g_sensor_int_s1_readdata;                           // g_sensor_int:readdata -> mm_interconnect_1:g_sensor_int_s1_readdata
	wire   [0:0] clock_crossing_io_m0_burstcount;                                      // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire         clock_crossing_io_m0_waitrequest;                                     // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire   [6:0] clock_crossing_io_m0_address;                                         // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire  [31:0] clock_crossing_io_m0_writedata;                                       // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                           // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire         clock_crossing_io_m0_read;                                            // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire  [31:0] clock_crossing_io_m0_readdata;                                        // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                                     // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire   [3:0] clock_crossing_io_m0_byteenable;                                      // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                                   // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire   [0:0] clock_crossing_io2_m0_burstcount;                                     // clock_crossing_io2:m0_burstcount -> mm_interconnect_2:clock_crossing_io2_m0_burstcount
	wire         clock_crossing_io2_m0_waitrequest;                                    // mm_interconnect_2:clock_crossing_io2_m0_waitrequest -> clock_crossing_io2:m0_waitrequest
	wire  [11:0] clock_crossing_io2_m0_address;                                        // clock_crossing_io2:m0_address -> mm_interconnect_2:clock_crossing_io2_m0_address
	wire  [31:0] clock_crossing_io2_m0_writedata;                                      // clock_crossing_io2:m0_writedata -> mm_interconnect_2:clock_crossing_io2_m0_writedata
	wire         clock_crossing_io2_m0_write;                                          // clock_crossing_io2:m0_write -> mm_interconnect_2:clock_crossing_io2_m0_write
	wire         clock_crossing_io2_m0_read;                                           // clock_crossing_io2:m0_read -> mm_interconnect_2:clock_crossing_io2_m0_read
	wire  [31:0] clock_crossing_io2_m0_readdata;                                       // mm_interconnect_2:clock_crossing_io2_m0_readdata -> clock_crossing_io2:m0_readdata
	wire         clock_crossing_io2_m0_debugaccess;                                    // clock_crossing_io2:m0_debugaccess -> mm_interconnect_2:clock_crossing_io2_m0_debugaccess
	wire   [3:0] clock_crossing_io2_m0_byteenable;                                     // clock_crossing_io2:m0_byteenable -> mm_interconnect_2:clock_crossing_io2_m0_byteenable
	wire         clock_crossing_io2_m0_readdatavalid;                                  // mm_interconnect_2:clock_crossing_io2_m0_readdatavalid -> clock_crossing_io2:m0_readdatavalid
	wire  [31:0] mm_interconnect_2_epcs_epcs_control_port_writedata;                   // mm_interconnect_2:epcs_epcs_control_port_writedata -> epcs:writedata
	wire   [8:0] mm_interconnect_2_epcs_epcs_control_port_address;                     // mm_interconnect_2:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_2_epcs_epcs_control_port_chipselect;                  // mm_interconnect_2:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire         mm_interconnect_2_epcs_epcs_control_port_write;                       // mm_interconnect_2:epcs_epcs_control_port_write -> epcs:write_n
	wire         mm_interconnect_2_epcs_epcs_control_port_read;                        // mm_interconnect_2:epcs_epcs_control_port_read -> epcs:read_n
	wire  [31:0] mm_interconnect_2_epcs_epcs_control_port_readdata;                    // epcs:readdata -> mm_interconnect_2:epcs_epcs_control_port_readdata
	wire   [7:0] mm_interconnect_2_gsensor_spi_slave_writedata;                        // mm_interconnect_2:gsensor_spi_slave_writedata -> gsensor_spi:s_writedata
	wire   [3:0] mm_interconnect_2_gsensor_spi_slave_address;                          // mm_interconnect_2:gsensor_spi_slave_address -> gsensor_spi:s_address
	wire         mm_interconnect_2_gsensor_spi_slave_chipselect;                       // mm_interconnect_2:gsensor_spi_slave_chipselect -> gsensor_spi:s_chipselect
	wire         mm_interconnect_2_gsensor_spi_slave_write;                            // mm_interconnect_2:gsensor_spi_slave_write -> gsensor_spi:s_write
	wire         mm_interconnect_2_gsensor_spi_slave_read;                             // mm_interconnect_2:gsensor_spi_slave_read -> gsensor_spi:s_read
	wire   [7:0] mm_interconnect_2_gsensor_spi_slave_readdata;                         // gsensor_spi:s_readdata -> mm_interconnect_2:gsensor_spi_slave_readdata
	wire  [31:0] mm_interconnect_2_i2c_scl_s1_writedata;                               // mm_interconnect_2:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire   [1:0] mm_interconnect_2_i2c_scl_s1_address;                                 // mm_interconnect_2:i2c_scl_s1_address -> i2c_scl:address
	wire         mm_interconnect_2_i2c_scl_s1_chipselect;                              // mm_interconnect_2:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire         mm_interconnect_2_i2c_scl_s1_write;                                   // mm_interconnect_2:i2c_scl_s1_write -> i2c_scl:write_n
	wire  [31:0] mm_interconnect_2_i2c_scl_s1_readdata;                                // i2c_scl:readdata -> mm_interconnect_2:i2c_scl_s1_readdata
	wire  [31:0] mm_interconnect_2_i2c_sda_s1_writedata;                               // mm_interconnect_2:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire   [1:0] mm_interconnect_2_i2c_sda_s1_address;                                 // mm_interconnect_2:i2c_sda_s1_address -> i2c_sda:address
	wire         mm_interconnect_2_i2c_sda_s1_chipselect;                              // mm_interconnect_2:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire         mm_interconnect_2_i2c_sda_s1_write;                                   // mm_interconnect_2:i2c_sda_s1_write -> i2c_sda:write_n
	wire  [31:0] mm_interconnect_2_i2c_sda_s1_readdata;                                // i2c_sda:readdata -> mm_interconnect_2:i2c_sda_s1_readdata
	wire         irq_mapper_receiver4_irq;                                             // jtag_uart:av_irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_d_irq_irq;                                                        // irq_mapper:sender_irq -> cpu:d_irq
	wire         irq_mapper_receiver0_irq;                                             // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                        // key:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                             // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                    // sw:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                             // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                    // g_sensor_int:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                             // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                                    // epcs:irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver5_irq;                                             // irq_synchronizer_004:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                                    // controller_interrupt_counter:irq -> irq_synchronizer_004:receiver_irq
	wire         irq_mapper_receiver6_irq;                                             // irq_synchronizer_005:sender_irq -> irq_mapper:receiver6_irq
	wire   [0:0] irq_synchronizer_005_receiver_irq;                                    // power_management_slave_0:error -> irq_synchronizer_005:receiver_irq
	wire         irq_mapper_receiver7_irq;                                             // irq_synchronizer_006:sender_irq -> irq_mapper:receiver7_irq
	wire   [0:0] irq_synchronizer_006_receiver_irq;                                    // RS232_0:irq -> irq_synchronizer_006:receiver_irq
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [clock_crossing_io:m0_reset, g_sensor_int:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, key:reset_n, led:reset_n, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset, select_i2c_clk:reset_n, sw:reset_n, sysid:reset_n]
	wire         cpu_jtag_debug_module_reset_reset;                                    // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [RS232_0:reset, altpll_sys:reset, clock_crossing_io2:m0_reset, controller_interrupt_counter:reset_n, epcs:reset_n, gsensor_spi:reset_n, i2c_scl:reset_n, i2c_sda:reset_n, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, mm_interconnect_0:altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset, mm_interconnect_2:clock_crossing_io2_m0_reset_reset_bridge_in_reset_reset, motor_controller_0:reset, power_management_slave_0:reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                               // rst_controller_001:reset_req -> [epcs:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                                   // rst_controller_002:reset_out -> [clock_crossing_io2:s0_reset, clock_crossing_io:s0_reset, cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_translator_001:in_reset, sdram:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                               // rst_controller_002:reset_req -> [cpu:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                                   // rst_controller_003:reset_out -> [imu_controller_0:spi_reset, mm_interconnect_0:imu_controller_0_reset_sink_reset_bridge_in_reset_reset]

	DE0_Nano_SOPC_key key (
		.clk        (altpll_io),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_key),                  // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)        //                 irq.irq
	);

	DE0_Nano_SOPC_sw sw (
		.clk        (altpll_io),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_sw),                  // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)   //                 irq.irq
	);

	DE0_Nano_SOPC_led led (
		.clk        (altpll_io),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led)                // external_connection.export
	);

	DE0_Nano_SOPC_i2c_scl i2c_scl (
		.clk        (clk_50),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_2_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_i2c_scl)                // external_connection.export
	);

	DE0_Nano_SOPC_i2c_sda i2c_sda (
		.clk        (clk_50),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_2_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (bidir_port_to_and_from_the_i2c_sda)       // external_connection.export
	);

	DE0_Nano_SOPC_sdram sdram (
		.clk            (altpll_sys),                               //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                   //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                     //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                  //      .export
		.zs_cke         (zs_cke_from_the_sdram),                    //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                   //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),              //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                    //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                  //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                    //      .export
	);

	DE0_Nano_SOPC_altpll_sys altpll_sys_inst (
		.clk       (clk_50),                                           //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),               // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_sys_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_sys_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_sys_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_sys_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_sys_pll_slave_writedata), //                      .writedata
		.c0        (altpll_sys),                                       //                    c0.clk
		.c1        (altpll_sdram),                                     //                    c1.clk
		.c2        (altpll_io),                                        //                    c2.clk
		.c3        (altpll_sys_c3_out),                                //                    c3.clk
		.c4        (altpll_adc),                                       //                    c4.clk
		.locked    (locked_from_the_altpll_sys),                       //        locked_conduit.export
		.phasedone (phasedone_from_the_altpll_sys)                     //     phasedone_conduit.export
	);

	DE0_Nano_SOPC_g_sensor_int g_sensor_int (
		.clk        (altpll_io),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_g_sensor_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_g_sensor_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_g_sensor_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_g_sensor_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_g_sensor_int_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_g_sensor_int),                  // external_connection.export
		.irq        (irq_synchronizer_002_receiver_irq)             //                 irq.irq
	);

	DE0_Nano_SOPC_epcs epcs (
		.clk           (clk_50),                                              //               clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                 //             reset.reset_n
		.reset_req     (rst_controller_001_reset_out_reset_req),              //                  .reset_req
		.address       (mm_interconnect_2_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_2_epcs_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                    //                  .dataavailable
		.endofpacket   (),                                                    //                  .endofpacket
		.read_n        (~mm_interconnect_2_epcs_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_2_epcs_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                    //                  .readyfordata
		.write_n       (~mm_interconnect_2_epcs_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_2_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_synchronizer_003_receiver_irq),                   //               irq.irq
		.dclk          (dclk_from_the_epcs),                                  //          external.export
		.sce           (sce_from_the_epcs),                                   //                  .export
		.sdo           (sdo_from_the_epcs),                                   //                  .export
		.data0         (data0_to_the_epcs)                                    //                  .export
	);

	DE0_Nano_SOPC_jtag_uart jtag_uart (
		.clk            (altpll_sys),                                                //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver4_irq)                                   //               irq.irq
	);

	TERASIC_SPI_3WIRE gsensor_spi (
		.clk          (clk_50),                                         //       clock_reset.clk
		.reset_n      (~rst_controller_001_reset_out_reset),            // clock_reset_reset.reset_n
		.s_chipselect (mm_interconnect_2_gsensor_spi_slave_chipselect), //             slave.chipselect
		.s_address    (mm_interconnect_2_gsensor_spi_slave_address),    //                  .address
		.s_write      (mm_interconnect_2_gsensor_spi_slave_write),      //                  .write
		.s_writedata  (mm_interconnect_2_gsensor_spi_slave_writedata),  //                  .writedata
		.s_read       (mm_interconnect_2_gsensor_spi_slave_read),       //                  .read
		.s_readdata   (mm_interconnect_2_gsensor_spi_slave_readdata),   //                  .readdata
		.SPI_SDIO     (SPI_SDIO_to_and_from_the_gsensor_spi),           //       conduit_end.export
		.SPI_SCLK     (SPI_SCLK_from_the_gsensor_spi),                  //                  .export
		.SPI_CS_n     (SPI_CS_n_from_the_gsensor_spi)                   //                  .export
	);

	DE0_Nano_SOPC_select_i2c_clk select_i2c_clk (
		.clk        (altpll_io),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_1_select_i2c_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_select_i2c_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_select_i2c_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_select_i2c_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_select_i2c_clk_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_select_i2c_clk)                // external_connection.export
	);

	slave_controller motor_controller_0 (
		.clk        (clk_50),                                                         //          clock.clk
		.chipselect (mm_interconnect_0_motor_controller_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.write      (mm_interconnect_0_motor_controller_0_avalon_slave_0_write),      //               .write
		.addr       (mm_interconnect_0_motor_controller_0_avalon_slave_0_address),    //               .address
		.writedata  (mm_interconnect_0_motor_controller_0_avalon_slave_0_writedata),  //               .writedata
		.GPIO_out   (GPIO_out_from_the_motor_controller_0),                           //    conduit_end.export
		.reset      (rst_controller_001_reset_out_reset)                              //          reset.reset
	);

	DE0_Nano_SOPC_controller_interrupt_counter controller_interrupt_counter (
		.clk        (clk_50),                                                       //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                          // reset.reset_n
		.address    (mm_interconnect_0_controller_interrupt_counter_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_controller_interrupt_counter_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_controller_interrupt_counter_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_controller_interrupt_counter_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_controller_interrupt_counter_s1_write),     //      .write_n
		.irq        (irq_synchronizer_004_receiver_irq)                             //   irq.irq
	);

	power_management_slave power_management_slave_0 (
		.chipselect (mm_interconnect_0_power_management_slave_0_avalon_slave_0_chipselect), //   avalon_slave_0.chipselect
		.write      (mm_interconnect_0_power_management_slave_0_avalon_slave_0_write),      //                 .write
		.read       (mm_interconnect_0_power_management_slave_0_avalon_slave_0_read),       //                 .read
		.writedata  (mm_interconnect_0_power_management_slave_0_avalon_slave_0_writedata),  //                 .writedata
		.readdata   (mm_interconnect_0_power_management_slave_0_avalon_slave_0_readdata),   //                 .readdata
		.clk        (clk_50),                                                               //            clock.clk
		.kill_sw    (kill_sw_from_the_power_management_slave_0),                            //      conduit_end.export
		.mux        (mux_from_the_power_management_slave_0),                                //                 .export
		.data       (data_to_the_power_management_slave_0),                                 //                 .export
		.error      (irq_synchronizer_005_receiver_irq),                                    // interrupt_sender.irq
		.reset      (rst_controller_001_reset_out_reset)                                    //            reset.reset
	);

	imu_controller imu_controller_0 (
		.spi_clk    (altpll_adc),                                                   //          clock.clk
		.chipselect (mm_interconnect_0_imu_controller_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.addr       (mm_interconnect_0_imu_controller_0_avalon_slave_0_address),    //               .address
		.read       (mm_interconnect_0_imu_controller_0_avalon_slave_0_read),       //               .read
		.readdata   (mm_interconnect_0_imu_controller_0_avalon_slave_0_readdata),   //               .readdata
		.sys_clk    (sys_clk_to_the_imu_controller_0),                              //    conduit_end.export
		.ADC_SDAT   (ADC_SDAT_to_the_imu_controller_0),                             //               .export
		.ADC_CS_N   (ADC_CS_N_from_the_imu_controller_0),                           //               .export
		.ADC_SADDR  (ADC_SADDR_from_the_imu_controller_0),                          //               .export
		.ADC_SCLK   (ADC_SCLK_from_the_imu_controller_0),                           //               .export
		.spi_reset  (rst_controller_003_reset_out_reset)                            //     reset_sink.reset
	);

	Altera_UP_Avalon_RS232 rs232_0 (
		.clk        (clk_50),                                              //            clock.clk
		.reset      (rst_controller_001_reset_out_reset),                  //            reset.reset
		.address    (mm_interconnect_0_rs232_0_avalon_slave_0_address),    //   avalon_slave_0.address
		.chipselect (mm_interconnect_0_rs232_0_avalon_slave_0_chipselect), //                 .chipselect
		.byteenable (mm_interconnect_0_rs232_0_avalon_slave_0_byteenable), //                 .byteenable
		.read       (mm_interconnect_0_rs232_0_avalon_slave_0_read),       //                 .read
		.write      (mm_interconnect_0_rs232_0_avalon_slave_0_write),      //                 .write
		.writedata  (mm_interconnect_0_rs232_0_avalon_slave_0_writedata),  //                 .writedata
		.readdata   (mm_interconnect_0_rs232_0_avalon_slave_0_readdata),   //                 .readdata
		.UART_RXD   (UART_RXD_to_the_RS232_0),                             //      conduit_end.export
		.UART_TXD   (UART_TXD_from_the_RS232_0),                           //    conduit_end_1.export
		.irq        (irq_synchronizer_006_receiver_irq)                    // interrupt_sender.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (7),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (altpll_io),                                            //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                       // m0_reset.reset
		.s0_clk           (altpll_sys),                                           //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (12),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io2 (
		.m0_clk           (clk_50),                                                //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                    // m0_reset.reset
		.s0_clk           (altpll_sys),                                            //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                    // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io2_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io2_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io2_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io2_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io2_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io2_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io2_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io2_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io2_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io2_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io2_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io2_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io2_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io2_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io2_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io2_m0_address),                         //         .address
		.m0_write         (clock_crossing_io2_m0_write),                           //         .write
		.m0_read          (clock_crossing_io2_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io2_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io2_m0_debugaccess)                      //         .debugaccess
	);

	DE0_Nano_SOPC_cpu cpu (
		.clk                                   (altpll_sys),                                          //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	DE0_Nano_SOPC_sysid sysid (
		.clock    (altpll_io),                                      //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	DE0_Nano_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.altpll_sys_c0_clk                                            (altpll_sys),                                                           //                                          altpll_sys_c0.clk
		.altpll_sys_c4_clk                                            (altpll_adc),                                                           //                                          altpll_sys_c4.clk
		.clk_50_clk_clk                                               (clk_50),                                                               //                                             clk_50_clk.clk
		.altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                   // altpll_sys_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_reset_n_reset_bridge_in_reset_reset                      (rst_controller_002_reset_out_reset),                                   //                      cpu_reset_n_reset_bridge_in_reset.reset
		.imu_controller_0_reset_sink_reset_bridge_in_reset_reset      (rst_controller_003_reset_out_reset),                                   //      imu_controller_0_reset_sink_reset_bridge_in_reset.reset
		.cpu_data_master_address                                      (cpu_data_master_address),                                              //                                        cpu_data_master.address
		.cpu_data_master_waitrequest                                  (cpu_data_master_waitrequest),                                          //                                                       .waitrequest
		.cpu_data_master_byteenable                                   (cpu_data_master_byteenable),                                           //                                                       .byteenable
		.cpu_data_master_read                                         (cpu_data_master_read),                                                 //                                                       .read
		.cpu_data_master_readdata                                     (cpu_data_master_readdata),                                             //                                                       .readdata
		.cpu_data_master_write                                        (cpu_data_master_write),                                                //                                                       .write
		.cpu_data_master_writedata                                    (cpu_data_master_writedata),                                            //                                                       .writedata
		.cpu_data_master_debugaccess                                  (cpu_data_master_debugaccess),                                          //                                                       .debugaccess
		.cpu_instruction_master_address                               (cpu_instruction_master_address),                                       //                                 cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                           (cpu_instruction_master_waitrequest),                                   //                                                       .waitrequest
		.cpu_instruction_master_read                                  (cpu_instruction_master_read),                                          //                                                       .read
		.cpu_instruction_master_readdata                              (cpu_instruction_master_readdata),                                      //                                                       .readdata
		.altpll_sys_pll_slave_address                                 (mm_interconnect_0_altpll_sys_pll_slave_address),                       //                                   altpll_sys_pll_slave.address
		.altpll_sys_pll_slave_write                                   (mm_interconnect_0_altpll_sys_pll_slave_write),                         //                                                       .write
		.altpll_sys_pll_slave_read                                    (mm_interconnect_0_altpll_sys_pll_slave_read),                          //                                                       .read
		.altpll_sys_pll_slave_readdata                                (mm_interconnect_0_altpll_sys_pll_slave_readdata),                      //                                                       .readdata
		.altpll_sys_pll_slave_writedata                               (mm_interconnect_0_altpll_sys_pll_slave_writedata),                     //                                                       .writedata
		.clock_crossing_io_s0_address                                 (mm_interconnect_0_clock_crossing_io_s0_address),                       //                                   clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                                   (mm_interconnect_0_clock_crossing_io_s0_write),                         //                                                       .write
		.clock_crossing_io_s0_read                                    (mm_interconnect_0_clock_crossing_io_s0_read),                          //                                                       .read
		.clock_crossing_io_s0_readdata                                (mm_interconnect_0_clock_crossing_io_s0_readdata),                      //                                                       .readdata
		.clock_crossing_io_s0_writedata                               (mm_interconnect_0_clock_crossing_io_s0_writedata),                     //                                                       .writedata
		.clock_crossing_io_s0_burstcount                              (mm_interconnect_0_clock_crossing_io_s0_burstcount),                    //                                                       .burstcount
		.clock_crossing_io_s0_byteenable                              (mm_interconnect_0_clock_crossing_io_s0_byteenable),                    //                                                       .byteenable
		.clock_crossing_io_s0_readdatavalid                           (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),                 //                                                       .readdatavalid
		.clock_crossing_io_s0_waitrequest                             (mm_interconnect_0_clock_crossing_io_s0_waitrequest),                   //                                                       .waitrequest
		.clock_crossing_io_s0_debugaccess                             (mm_interconnect_0_clock_crossing_io_s0_debugaccess),                   //                                                       .debugaccess
		.clock_crossing_io2_s0_address                                (mm_interconnect_0_clock_crossing_io2_s0_address),                      //                                  clock_crossing_io2_s0.address
		.clock_crossing_io2_s0_write                                  (mm_interconnect_0_clock_crossing_io2_s0_write),                        //                                                       .write
		.clock_crossing_io2_s0_read                                   (mm_interconnect_0_clock_crossing_io2_s0_read),                         //                                                       .read
		.clock_crossing_io2_s0_readdata                               (mm_interconnect_0_clock_crossing_io2_s0_readdata),                     //                                                       .readdata
		.clock_crossing_io2_s0_writedata                              (mm_interconnect_0_clock_crossing_io2_s0_writedata),                    //                                                       .writedata
		.clock_crossing_io2_s0_burstcount                             (mm_interconnect_0_clock_crossing_io2_s0_burstcount),                   //                                                       .burstcount
		.clock_crossing_io2_s0_byteenable                             (mm_interconnect_0_clock_crossing_io2_s0_byteenable),                   //                                                       .byteenable
		.clock_crossing_io2_s0_readdatavalid                          (mm_interconnect_0_clock_crossing_io2_s0_readdatavalid),                //                                                       .readdatavalid
		.clock_crossing_io2_s0_waitrequest                            (mm_interconnect_0_clock_crossing_io2_s0_waitrequest),                  //                                                       .waitrequest
		.clock_crossing_io2_s0_debugaccess                            (mm_interconnect_0_clock_crossing_io2_s0_debugaccess),                  //                                                       .debugaccess
		.controller_interrupt_counter_s1_address                      (mm_interconnect_0_controller_interrupt_counter_s1_address),            //                        controller_interrupt_counter_s1.address
		.controller_interrupt_counter_s1_write                        (mm_interconnect_0_controller_interrupt_counter_s1_write),              //                                                       .write
		.controller_interrupt_counter_s1_readdata                     (mm_interconnect_0_controller_interrupt_counter_s1_readdata),           //                                                       .readdata
		.controller_interrupt_counter_s1_writedata                    (mm_interconnect_0_controller_interrupt_counter_s1_writedata),          //                                                       .writedata
		.controller_interrupt_counter_s1_chipselect                   (mm_interconnect_0_controller_interrupt_counter_s1_chipselect),         //                                                       .chipselect
		.cpu_jtag_debug_module_address                                (mm_interconnect_0_cpu_jtag_debug_module_address),                      //                                  cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                                  (mm_interconnect_0_cpu_jtag_debug_module_write),                        //                                                       .write
		.cpu_jtag_debug_module_read                                   (mm_interconnect_0_cpu_jtag_debug_module_read),                         //                                                       .read
		.cpu_jtag_debug_module_readdata                               (mm_interconnect_0_cpu_jtag_debug_module_readdata),                     //                                                       .readdata
		.cpu_jtag_debug_module_writedata                              (mm_interconnect_0_cpu_jtag_debug_module_writedata),                    //                                                       .writedata
		.cpu_jtag_debug_module_byteenable                             (mm_interconnect_0_cpu_jtag_debug_module_byteenable),                   //                                                       .byteenable
		.cpu_jtag_debug_module_waitrequest                            (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),                  //                                                       .waitrequest
		.cpu_jtag_debug_module_debugaccess                            (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),                  //                                                       .debugaccess
		.imu_controller_0_avalon_slave_0_address                      (mm_interconnect_0_imu_controller_0_avalon_slave_0_address),            //                        imu_controller_0_avalon_slave_0.address
		.imu_controller_0_avalon_slave_0_read                         (mm_interconnect_0_imu_controller_0_avalon_slave_0_read),               //                                                       .read
		.imu_controller_0_avalon_slave_0_readdata                     (mm_interconnect_0_imu_controller_0_avalon_slave_0_readdata),           //                                                       .readdata
		.imu_controller_0_avalon_slave_0_chipselect                   (mm_interconnect_0_imu_controller_0_avalon_slave_0_chipselect),         //                                                       .chipselect
		.jtag_uart_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                //                            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                  //                                                       .write
		.jtag_uart_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                   //                                                       .read
		.jtag_uart_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),               //                                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),              //                                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),            //                                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),             //                                                       .chipselect
		.motor_controller_0_avalon_slave_0_address                    (mm_interconnect_0_motor_controller_0_avalon_slave_0_address),          //                      motor_controller_0_avalon_slave_0.address
		.motor_controller_0_avalon_slave_0_write                      (mm_interconnect_0_motor_controller_0_avalon_slave_0_write),            //                                                       .write
		.motor_controller_0_avalon_slave_0_writedata                  (mm_interconnect_0_motor_controller_0_avalon_slave_0_writedata),        //                                                       .writedata
		.motor_controller_0_avalon_slave_0_chipselect                 (mm_interconnect_0_motor_controller_0_avalon_slave_0_chipselect),       //                                                       .chipselect
		.power_management_slave_0_avalon_slave_0_write                (mm_interconnect_0_power_management_slave_0_avalon_slave_0_write),      //                power_management_slave_0_avalon_slave_0.write
		.power_management_slave_0_avalon_slave_0_read                 (mm_interconnect_0_power_management_slave_0_avalon_slave_0_read),       //                                                       .read
		.power_management_slave_0_avalon_slave_0_readdata             (mm_interconnect_0_power_management_slave_0_avalon_slave_0_readdata),   //                                                       .readdata
		.power_management_slave_0_avalon_slave_0_writedata            (mm_interconnect_0_power_management_slave_0_avalon_slave_0_writedata),  //                                                       .writedata
		.power_management_slave_0_avalon_slave_0_chipselect           (mm_interconnect_0_power_management_slave_0_avalon_slave_0_chipselect), //                                                       .chipselect
		.RS232_0_avalon_slave_0_address                               (mm_interconnect_0_rs232_0_avalon_slave_0_address),                     //                                 RS232_0_avalon_slave_0.address
		.RS232_0_avalon_slave_0_write                                 (mm_interconnect_0_rs232_0_avalon_slave_0_write),                       //                                                       .write
		.RS232_0_avalon_slave_0_read                                  (mm_interconnect_0_rs232_0_avalon_slave_0_read),                        //                                                       .read
		.RS232_0_avalon_slave_0_readdata                              (mm_interconnect_0_rs232_0_avalon_slave_0_readdata),                    //                                                       .readdata
		.RS232_0_avalon_slave_0_writedata                             (mm_interconnect_0_rs232_0_avalon_slave_0_writedata),                   //                                                       .writedata
		.RS232_0_avalon_slave_0_byteenable                            (mm_interconnect_0_rs232_0_avalon_slave_0_byteenable),                  //                                                       .byteenable
		.RS232_0_avalon_slave_0_chipselect                            (mm_interconnect_0_rs232_0_avalon_slave_0_chipselect),                  //                                                       .chipselect
		.sdram_s1_address                                             (mm_interconnect_0_sdram_s1_address),                                   //                                               sdram_s1.address
		.sdram_s1_write                                               (mm_interconnect_0_sdram_s1_write),                                     //                                                       .write
		.sdram_s1_read                                                (mm_interconnect_0_sdram_s1_read),                                      //                                                       .read
		.sdram_s1_readdata                                            (mm_interconnect_0_sdram_s1_readdata),                                  //                                                       .readdata
		.sdram_s1_writedata                                           (mm_interconnect_0_sdram_s1_writedata),                                 //                                                       .writedata
		.sdram_s1_byteenable                                          (mm_interconnect_0_sdram_s1_byteenable),                                //                                                       .byteenable
		.sdram_s1_readdatavalid                                       (mm_interconnect_0_sdram_s1_readdatavalid),                             //                                                       .readdatavalid
		.sdram_s1_waitrequest                                         (mm_interconnect_0_sdram_s1_waitrequest),                               //                                                       .waitrequest
		.sdram_s1_chipselect                                          (mm_interconnect_0_sdram_s1_chipselect)                                 //                                                       .chipselect
	);

	DE0_Nano_SOPC_mm_interconnect_1 mm_interconnect_1 (
		.altpll_sys_c2_clk                                      (altpll_io),                                      //                                    altpll_sys_c2.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                 // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                   //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),               //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                      //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                  //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),             //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                     //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                 //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),               //                                                 .debugaccess
		.g_sensor_int_s1_address                                (mm_interconnect_1_g_sensor_int_s1_address),      //                                  g_sensor_int_s1.address
		.g_sensor_int_s1_write                                  (mm_interconnect_1_g_sensor_int_s1_write),        //                                                 .write
		.g_sensor_int_s1_readdata                               (mm_interconnect_1_g_sensor_int_s1_readdata),     //                                                 .readdata
		.g_sensor_int_s1_writedata                              (mm_interconnect_1_g_sensor_int_s1_writedata),    //                                                 .writedata
		.g_sensor_int_s1_chipselect                             (mm_interconnect_1_g_sensor_int_s1_chipselect),   //                                                 .chipselect
		.key_s1_address                                         (mm_interconnect_1_key_s1_address),               //                                           key_s1.address
		.key_s1_write                                           (mm_interconnect_1_key_s1_write),                 //                                                 .write
		.key_s1_readdata                                        (mm_interconnect_1_key_s1_readdata),              //                                                 .readdata
		.key_s1_writedata                                       (mm_interconnect_1_key_s1_writedata),             //                                                 .writedata
		.key_s1_chipselect                                      (mm_interconnect_1_key_s1_chipselect),            //                                                 .chipselect
		.led_s1_address                                         (mm_interconnect_1_led_s1_address),               //                                           led_s1.address
		.led_s1_write                                           (mm_interconnect_1_led_s1_write),                 //                                                 .write
		.led_s1_readdata                                        (mm_interconnect_1_led_s1_readdata),              //                                                 .readdata
		.led_s1_writedata                                       (mm_interconnect_1_led_s1_writedata),             //                                                 .writedata
		.led_s1_chipselect                                      (mm_interconnect_1_led_s1_chipselect),            //                                                 .chipselect
		.select_i2c_clk_s1_address                              (mm_interconnect_1_select_i2c_clk_s1_address),    //                                select_i2c_clk_s1.address
		.select_i2c_clk_s1_write                                (mm_interconnect_1_select_i2c_clk_s1_write),      //                                                 .write
		.select_i2c_clk_s1_readdata                             (mm_interconnect_1_select_i2c_clk_s1_readdata),   //                                                 .readdata
		.select_i2c_clk_s1_writedata                            (mm_interconnect_1_select_i2c_clk_s1_writedata),  //                                                 .writedata
		.select_i2c_clk_s1_chipselect                           (mm_interconnect_1_select_i2c_clk_s1_chipselect), //                                                 .chipselect
		.sw_s1_address                                          (mm_interconnect_1_sw_s1_address),                //                                            sw_s1.address
		.sw_s1_write                                            (mm_interconnect_1_sw_s1_write),                  //                                                 .write
		.sw_s1_readdata                                         (mm_interconnect_1_sw_s1_readdata),               //                                                 .readdata
		.sw_s1_writedata                                        (mm_interconnect_1_sw_s1_writedata),              //                                                 .writedata
		.sw_s1_chipselect                                       (mm_interconnect_1_sw_s1_chipselect),             //                                                 .chipselect
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),  //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata)  //                                                 .readdata
	);

	DE0_Nano_SOPC_mm_interconnect_2 mm_interconnect_2 (
		.clk_50_clk_clk                                          (clk_50),                                              //                                        clk_50_clk.clk
		.clock_crossing_io2_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                  // clock_crossing_io2_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_io2_m0_address                           (clock_crossing_io2_m0_address),                       //                             clock_crossing_io2_m0.address
		.clock_crossing_io2_m0_waitrequest                       (clock_crossing_io2_m0_waitrequest),                   //                                                  .waitrequest
		.clock_crossing_io2_m0_burstcount                        (clock_crossing_io2_m0_burstcount),                    //                                                  .burstcount
		.clock_crossing_io2_m0_byteenable                        (clock_crossing_io2_m0_byteenable),                    //                                                  .byteenable
		.clock_crossing_io2_m0_read                              (clock_crossing_io2_m0_read),                          //                                                  .read
		.clock_crossing_io2_m0_readdata                          (clock_crossing_io2_m0_readdata),                      //                                                  .readdata
		.clock_crossing_io2_m0_readdatavalid                     (clock_crossing_io2_m0_readdatavalid),                 //                                                  .readdatavalid
		.clock_crossing_io2_m0_write                             (clock_crossing_io2_m0_write),                         //                                                  .write
		.clock_crossing_io2_m0_writedata                         (clock_crossing_io2_m0_writedata),                     //                                                  .writedata
		.clock_crossing_io2_m0_debugaccess                       (clock_crossing_io2_m0_debugaccess),                   //                                                  .debugaccess
		.epcs_epcs_control_port_address                          (mm_interconnect_2_epcs_epcs_control_port_address),    //                            epcs_epcs_control_port.address
		.epcs_epcs_control_port_write                            (mm_interconnect_2_epcs_epcs_control_port_write),      //                                                  .write
		.epcs_epcs_control_port_read                             (mm_interconnect_2_epcs_epcs_control_port_read),       //                                                  .read
		.epcs_epcs_control_port_readdata                         (mm_interconnect_2_epcs_epcs_control_port_readdata),   //                                                  .readdata
		.epcs_epcs_control_port_writedata                        (mm_interconnect_2_epcs_epcs_control_port_writedata),  //                                                  .writedata
		.epcs_epcs_control_port_chipselect                       (mm_interconnect_2_epcs_epcs_control_port_chipselect), //                                                  .chipselect
		.gsensor_spi_slave_address                               (mm_interconnect_2_gsensor_spi_slave_address),         //                                 gsensor_spi_slave.address
		.gsensor_spi_slave_write                                 (mm_interconnect_2_gsensor_spi_slave_write),           //                                                  .write
		.gsensor_spi_slave_read                                  (mm_interconnect_2_gsensor_spi_slave_read),            //                                                  .read
		.gsensor_spi_slave_readdata                              (mm_interconnect_2_gsensor_spi_slave_readdata),        //                                                  .readdata
		.gsensor_spi_slave_writedata                             (mm_interconnect_2_gsensor_spi_slave_writedata),       //                                                  .writedata
		.gsensor_spi_slave_chipselect                            (mm_interconnect_2_gsensor_spi_slave_chipselect),      //                                                  .chipselect
		.i2c_scl_s1_address                                      (mm_interconnect_2_i2c_scl_s1_address),                //                                        i2c_scl_s1.address
		.i2c_scl_s1_write                                        (mm_interconnect_2_i2c_scl_s1_write),                  //                                                  .write
		.i2c_scl_s1_readdata                                     (mm_interconnect_2_i2c_scl_s1_readdata),               //                                                  .readdata
		.i2c_scl_s1_writedata                                    (mm_interconnect_2_i2c_scl_s1_writedata),              //                                                  .writedata
		.i2c_scl_s1_chipselect                                   (mm_interconnect_2_i2c_scl_s1_chipselect),             //                                                  .chipselect
		.i2c_sda_s1_address                                      (mm_interconnect_2_i2c_sda_s1_address),                //                                        i2c_sda_s1.address
		.i2c_sda_s1_write                                        (mm_interconnect_2_i2c_sda_s1_write),                  //                                                  .write
		.i2c_sda_s1_readdata                                     (mm_interconnect_2_i2c_sda_s1_readdata),               //                                                  .readdata
		.i2c_sda_s1_writedata                                    (mm_interconnect_2_i2c_sda_s1_writedata),              //                                                  .writedata
		.i2c_sda_s1_chipselect                                   (mm_interconnect_2_i2c_sda_s1_chipselect)              //                                                  .chipselect
	);

	DE0_Nano_SOPC_irq_mapper irq_mapper (
		.clk           (altpll_sys),                         //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),           // receiver7.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_io),                          //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_io),                          //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (altpll_io),                          //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_006 (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_006_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                          // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (altpll_io),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (clk_50),                                 //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (altpll_sys),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (altpll_adc),                         //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
